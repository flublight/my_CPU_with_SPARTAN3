`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/03/19 16:10:43
// Design Name:
// Module Name: IF_sim
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

`define WORD 32  // 1word
`define WORD_ADDR_W 30  // address width 1word

`define WORD_MSB `WORD-1
`define WORD_ADDR_MSB `WORD_ADDR_W-1


module IF_sim();
	reg				   clk=0;			// ????N????????????b????N
	reg				   reset;		// ???????????????????????????Z????b????g
	/********** SPM????C????????????^????t????F????[????X **********/
	reg [`WORD_MSB:0] spm_rd_data; // ????????�o????????????f????[????^
	wire [`WORD_ADDR_MSB:0] spm_addr;	// ????A????h????????????X
	wire				   spm_as_;		// ????A????h????????????X????X????g????????????[????u
	wire				   spm_rw;		// ?????????????????????????
	wire [`WORD_MSB:0] spm_wr_data; // ??????????????????????????????�R??[????^
	/********** ????o????X????C????????????^????t????F????[????X **********/
	reg [`WORD_MSB:0] bus_rd_data; // ????????�o????????????f????[????^
	reg				   bus_rdy_;	// ????????????f????B
	reg				   bus_grnt_;	// ????o????X????O????????????????????g
	wire				   bus_req_;	// ????o????X????????????N????G????X????g
	wire [`WORD_ADDR_MSB:0] bus_addr;	// ????A????h????????????X
	wire				   bus_as_;		// ????A????h????????????X????X????g????????????[????u
	wire				   bus_rw;		// ?????????????????????????
	wire [`WORD_MSB:0] bus_wr_data; // ??????????????????????????????�R??[????^
	/********** ????p????C????v????????????C????????????????????????????M???????? **********/
	reg				   stall;		// ????X????g????[????????
	reg				   flush;		// ????t????????????b????V????????
	reg [`WORD_ADDR_MSB:0] new_pc;		// ????V????????????????????v????????????O????????????????????J????E????????????^
	reg				   br_taken;	// ??????????????????????��????????????
	reg [`WORD_ADDR_MSB:0] br_addr;		// ????????????????????????????A????h????????????X
	wire				   busy;		// ????r????W????[????M????????
	/********** IF/ID????p????C????v????????????C????????????????????W????X????^ **********/
	wire [`WORD_ADDR_MSB:0] if_pc;		// ????v????????????O????????????????????J????E????????????^
	wire [`WORD_MSB:0] if_insn;		// ????????????????
	wire				   if_en;		// ????p????C????v????????????C????????????f????[????^??????��??????

	/********** ?????????????????????????????M???????? **********/
	wire [31:0]		   insn;		// ????t????F????b????`????????????????????????????????

	/********** ????o????X????C????????????^????t????F????[????X **********/
	bus_IF bus_if (
		/********** ????N????????????b????N & ????????????Z????b????g **********/
		.clk		 (clk),					// ????N????????????b????N
		.rst		 (reset),				// ???????????????????????????Z????b????g
		/********** ????p????C????v????????????C????????????????????????????M???????? **********/
		.stall		 (stall),				// ????X????g????[????????
		.flush		 (flush),				// ????t????????????b????V????????????M????????
		.busy		 (busy),				// ????r????W????[????M????????
		/********** CPU????C????????????^????t????F????[????X **********/
		.addr		 (if_pc),				// ????A????h????????????X
		.as		 (1'b1),			// ????A????h????????????X????L????????
		.rw			 (1'b0),				// ?????????????????????????
		.wr_data	 (32'h00000000),		// ??????????????????????????????�R??[????^
		.rd_data	 (insn),				// ????????�o????????????f????[????^
		/********** ????X????N????????????b????`????p????b????h????????????????????????????C????????????^????t????F????[????X **********/
		.spm_rd_data (spm_rd_data),			// ????????�o????????????f????[????^
		.spm_addr	 (spm_addr),			// ????A????h????????????X
		.spm_as	 (spm_as_),				// ????A????h????????????X????X????g????????????[????u
		.spm_rw		 (spm_rw),				// ?????????????????????????
		.spm_wr_data (spm_wr_data),			// ??????????????????????????????�R??[????^
		/********** ????o????X????C????????????^????t????F????[????X **********/
		.bus_rd_data (bus_rd_data),			// ????????�o????????????f????[????^
		.bus_rdy	 (bus_rdy_),			// ????????????f????B
		.bus_grnt	 (bus_grnt_),			// ????o????X????O????????????????????g
		.bus_req	 (bus_req_),			// ????o????X????????????N????G????X????g
		.bus_addr	 (bus_addr),			// ????A????h????????????X
		.bus_as	 (bus_as_),				// ????A????h????????????X????X????g????????????[????u
		.bus_rw		 (bus_rw),				// ?????????????????????????
		.bus_wr_data (bus_wr_data)			// ??????????????????????????????�R??[????^
	);

	/********** IF????X????e????[????W????p????C????v????????????C????????????????????W????X????^ **********/
	reg_IF if_reg (
		/********** ????N????????????b????N & ????????????Z????b????g **********/
		.clk		 (clk),					// ????N????????????b????N
		.rst		 (reset),				// ???????????????????????????Z????b????g
		/********** ????t????F????b????`????f????[????^ **********/
		.inst		 (insn),				// ????t????F????b????`????????????????????????????????
		/********** ????p????C????v????????????C????????????????????????????M???????? **********/
		.stall		 (stall),				// ????X????g????[????????
		.flush		 (flush),				// ????t????????????b????V????????
		.new_pc		 (new_pc),				// ????V????????????????????v????????????O????????????????????J????E????????????^
		.br_taken	 (br_taken),			// ??????????????????????��????????????
		.br_addr	 (br_addr),				// ????????????????????????????A????h????????????X
		/********** IF/ID????p????C????v????????????C????????????????????W????X????^ **********/
		.if_pc		 (if_pc),				// ????v????????????O????????????????????J????E????????????^
		.if_inst	 (if_insn),				// ????????????????
		.if_en		 (if_en)				// ????p????C????v????????????C????????????f????[????^??????��??????
	);


    always begin
       clk=~clk; #(5);
    end


  initial begin
    reset = 1;
		#(2)
    reset <= 0;
		repeat(2) @(posedge clk);
    reset <= 1;
		spm_rd_data=32'h00000001;
		bus_rd_data=32'h00000002; // ????????�o????????????f????[????^
		bus_rdy_=1;	// ????????????f????B
		bus_grnt_=1;	// ????o????X????O????????????????????g
		new_pc=30'h00001000;		//

		stall=0;
		flush=0;
    repeat(200) @(posedge clk);
		stall=0;
		flush=1;
    repeat(200) @(posedge clk);
		stall=1;
		flush=0;
    repeat(200) @(posedge clk);
		stall=1;
		flush=1;
		repeat(200) @(posedge clk);
		br_taken=0;	// ??????????????????????��????????????
		br_addr=30'h1000000;		// ????????????????????????????A????h????????????X
		stall=0;
		flush=0;
		repeat(200) @(posedge clk);

    $finish;
  end

endmodule
