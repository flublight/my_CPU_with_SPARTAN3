`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/03/07 16:35:44
// Design Name:
// Module Name: bus_IF
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

`define WORD 32  // 1word
`define WORD_ADDR_W 30  // address width 1word

`define WORD_MSB `WORD-1
`define WORD_ADDR_MSB `WORD_ADDR_W-1

module reg_IF (
  input clk,
  input rst,
  input[`WORD_MSB:0] inst,//fetch data(instraction)

  input stall,
  input flush,
  input[`WORD_ADDR_MSB:0] new_pc,
  input br_taken,
  input[`WORD_ADDR_MSB:0] br_addr,

  output reg[`WORD_ADDR_MSB:0] if_pc,
  output reg[`WORD_MSB:0] if_inst,
  output reg if_en
  );


  always@(posedge clk or negedge rst)begin//bus access control
    if(~rst)begin
      if_pc<=new_pc;
      if_inst<=0;//NOP
      if_en<=0;
    end
    else begin
      if(~stall)begin
        if(flush)begin
        if_pc<=new_pc;
        if_inst<=0;//NOP
        if_en<=0;
        end
        else if(br_taken)begin//branch
        if_pc<=br_addr;
        if_inst<=inst;//
        if_en<=1;
        end
        else begin
        if_pc<=if_pc+1;
        if_inst<=inst;//
        if_en<=1;
        end
      end
    end
 end
endmodule //if_reg

module bus_IF(
    input clk,
    input rst,
    input stall,
    input flush,
    output reg busy,
    //cpu_interface
    input [`WORD_ADDR_MSB:0]addr,
    input as,
    input rw,
    output reg [`WORD_MSB:0]rd_data,
    input [`WORD_MSB:0]wr_data,
    //spm
    input [`WORD_MSB:0]spm_rd_data,
    output [`WORD_ADDR_MSB:0]spm_addr,
    output reg spm_as,
    output spm_rw,
    output [`WORD_MSB:0]spm_wr_data,
    //bus
    input [`WORD_MSB:0]bus_rd_data,
    input bus_rdy,
    input bus_grnt,
    output reg[`WORD_ADDR_MSB:0]bus_addr,
    output reg[`WORD_MSB:0]bus_wr_data,
    output reg bus_req,
    output reg bus_rw,
    output reg bus_as
    );
reg [1:0]state;//0:idle,1:bus_req,2:bus_access,3:stull
reg[`WORD_MSB:0]rd_buf;
wire s_index;
assign s_index = addr[29:27];//slave_index

assign spm_rw=rw;
assign spm_wr_data=wr_data;
assign spm_addr=addr;



always@(*)begin//memory access control
      rd_data=0;
      spm_as=0;
      busy=0;
      case(state)
      0:begin
        if(~flush&&as)
          if(s_index==1)begin
            if(~stall)begin
              spm_as=1;
              if(rw==0)rd_data=spm_rd_data;//read
            end
          end
          else busy=1;
        end

      1:busy=1;

      2:begin
        if(bus_rdy)begin
          if(rw==0)rd_data=bus_rd_data;//read
        end
        else busy=1;
        end

      3:if(rw==0)rd_data=rd_buf;

      endcase
    end
    always@(posedge clk or negedge rst)begin//bus access control
      if(~rst)begin
        state<=0;
        bus_req<=0;
        bus_addr<=0;
        bus_as<=0;
        bus_rw<=0;
        bus_wr_data<=0;
        rd_buf<=0;
      end
      else begin
          case (state)
          0:
          if(~flush&&as)
            if(s_index!=1)begin
              state<=1;
              bus_req<=1;
              bus_addr<=addr;
              bus_rw<=rw;
              bus_wr_data<=wr_data;
          end
            1:if(bus_grnt)begin
                state<=2;
                bus_as<=1;
              end
            2:begin
                bus_as<=0;
                if(bus_rdy)begin
                bus_req<=0;
                bus_addr<=0;
                bus_rw<=0;
                bus_wr_data<=0;
                //store read data
                if(bus_rw==0)rd_buf<=bus_rd_data;

                //check stall
                if(stall)state<=3;
                else state<=0;
                end
              end

            3:if(~stall)state<=0;
          endcase
        end
     end
endmodule


module stage_IF (
	/********** ?�?�N?�?�?�?�?�?�b?�?�N & ?�?�?�?�?�?�Z?�?�b?�?�g **********/
	input  wire				   clk,			// ?�?�N?�?�?�?�?�?�b?�?�N
	input  wire				   reset,		// ?�?�������?��?�?�?�?�?�?�?�Z?�?�b?�?�g
	/********** SPM?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
	input  wire [`WORD_MSB:0] spm_rd_data, // ?�?�??��出?�?�?�?�?�?�f?�?�[?�?�^
	output wire [`WORD_ADDR_MSB:0] spm_addr,	// ?�?�A?�?�h?�?�?�?�?�?�X
	output wire				   spm_as_,		// ?�?�A?�?�h?�?�?�?�?�?�X?�?�X?�?�g?�?�?�?�?�?�[?�?�u
	output wire				   spm_rw,		// ?�?�??��?��?�?�?�?�?�?�?�
	output wire [`WORD_MSB:0] spm_wr_data, // ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�ヽ?�[?�?�^
	/********** ?�?�o?�?�X?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
	input  wire [`WORD_MSB:0] bus_rd_data, // ?�?�??��出?�?�?�?�?�?�f?�?�[?�?�^
	input  wire				   bus_rdy_,	// ?�?�?�?�?�?�f?�?�B
	input  wire				   bus_grnt_,	// ?�?�o?�?�X?�?�O?�?�?�?�?�?�?�?�?�?�g
	output wire				   bus_req_,	// ?�?�o?�?�X?�?�?�?�?�?�N?�?�G?�?�X?�?�g
	output wire [`WORD_ADDR_MSB:0] bus_addr,	// ?�?�A?�?�h?�?�?�?�?�?�X
	output wire				   bus_as_,		// ?�?�A?�?�h?�?�?�?�?�?�X?�?�X?�?�g?�?�?�?�?�?�[?�?�u
	output wire				   bus_rw,		// ?�?�??��?��?�?�?�?�?�?�?�
	output wire [`WORD_MSB:0] bus_wr_data, // ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�ヽ?�[?�?�^
	/********** ?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�?�?�?�?�M?�?�?�?� **********/
	input  wire				   stall,		// ?�?�X?�?�g?�?�[?�?�?�?�
	input  wire				   flush,		// ?�?�t?�?�?�?�?�?�b?�?�V?�?�?�?�
	input  wire [`WORD_ADDR_MSB:0] new_pc,		// ?�?�V?�?�?�?�?�?�?�?�?�?�v?�?�?�?�?�?�O?�?�?�?�?�?�?�?�?�?�J?�?�E?�?�?�?�?�?�^
	input  wire				   br_taken,	// ?�?�?�?�?�?�?�?�?�?�?�撰?�?�?�?�?�?�
	input  wire [`WORD_ADDR_MSB:0] br_addr,		// ?�?�?�?�?�?�?�?�?�?�?�?�?�?�A?�?�h?�?�?�?�?�?�X
	output wire				   busy,		// ?�?�r?�?�W?�?�[?�?�M?�?�?�?�
	/********** IF/ID?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�W?�?�X?�?�^ **********/
	output wire [`WORD_ADDR_MSB:0] if_pc,		// ?�?�v?�?�?�?�?�?�O?�?�?�?�?�?�?�?�?�?�J?�?�E?�?�?�?�?�?�^
	output wire [`WORD_MSB:0] if_insn,		// ?�?�?�?�?�?�?�?�
	output wire				   if_en		// ?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�f?�?�[?�?�^?�?�?�朽?�?�?�
);

	/********** ?�?�?�?�?�?�?�?�?�?�?�扽?�?�?�M?�?�?�?� **********/
	wire [31:0]		   insn;		// ?�?�t?�?�F?�?�b?�?�`?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�

	/********** ?�?�o?�?�X?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
	bus_IF bus_if (
		/********** ?�?�N?�?�?�?�?�?�b?�?�N & ?�?�?�?�?�?�Z?�?�b?�?�g **********/
		.clk		 (clk),					// ?�?�N?�?�?�?�?�?�b?�?�N
		.rst		 (reset),				// ?�?�������?��?�?�?�?�?�?�?�Z?�?�b?�?�g
		/********** ?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�?�?�?�?�M?�?�?�?� **********/
		.stall		 (stall),				// ?�?�X?�?�g?�?�[?�?�?�?�
		.flush		 (flush),				// ?�?�t?�?�?�?�?�?�b?�?�V?�?�?�?�?�?�M?�?�?�?�
		.busy		 (busy),				// ?�?�r?�?�W?�?�[?�?�M?�?�?�?�
		/********** CPU?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
		.addr		 (if_pc),				// ?�?�A?�?�h?�?�?�?�?�?�X
		.as		 (1'b1),			// ?�?�A?�?�h?�?�?�?�?�?�X?�?�L?�?�?�?�
		.rw			 (1'b0),				// ?�?�??��?��?�?�?�?�?�?�?�
		.wr_data	 (32'h00000000),		// ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�ヽ?�[?�?�^
		.rd_data	 (insn),				// ?�?�??��出?�?�?�?�?�?�f?�?�[?�?�^
		/********** ?�?�X?�?�N?�?�?�?�?�?�b?�?�`?�?�p?�?�b?�?�h?�?�?�?�?�?�?�?�?�?�?�?�?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
		.spm_rd_data (spm_rd_data),			// ?�?�??��出?�?�?�?�?�?�f?�?�[?�?�^
		.spm_addr	 (spm_addr),			// ?�?�A?�?�h?�?�?�?�?�?�X
		.spm_as	 (spm_as_),				// ?�?�A?�?�h?�?�?�?�?�?�X?�?�X?�?�g?�?�?�?�?�?�[?�?�u
		.spm_rw		 (spm_rw),				// ?�?�??��?��?�?�?�?�?�?�?�
		.spm_wr_data (spm_wr_data),			// ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�ヽ?�[?�?�^
		/********** ?�?�o?�?�X?�?�C?�?�?�?�?�?�^?�?�t?�?�F?�?�[?�?�X **********/
		.bus_rd_data (bus_rd_data),			// ?�?�??��出?�?�?�?�?�?�f?�?�[?�?�^
		.bus_rdy	 (bus_rdy_),			// ?�?�?�?�?�?�f?�?�B
		.bus_grnt	 (bus_grnt_),			// ?�?�o?�?�X?�?�O?�?�?�?�?�?�?�?�?�?�g
		.bus_req	 (bus_req_),			// ?�?�o?�?�X?�?�?�?�?�?�N?�?�G?�?�X?�?�g
		.bus_addr	 (bus_addr),			// ?�?�A?�?�h?�?�?�?�?�?�X
		.bus_as	 (bus_as_),				// ?�?�A?�?�h?�?�?�?�?�?�X?�?�X?�?�g?�?�?�?�?�?�[?�?�u
		.bus_rw		 (bus_rw),				// ?�?�??��?��?�?�?�?�?�?�?�
		.bus_wr_data (bus_wr_data)			// ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�ヽ?�[?�?�^
	);

	/********** IF?�?�X?�?�e?�?�[?�?�W?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�W?�?�X?�?�^ **********/
	reg_IF if_reg (
		/********** ?�?�N?�?�?�?�?�?�b?�?�N & ?�?�?�?�?�?�Z?�?�b?�?�g **********/
		.clk		 (clk),					// ?�?�N?�?�?�?�?�?�b?�?�N
		.rst		 (reset),				// ?�?�������?��?�?�?�?�?�?�?�Z?�?�b?�?�g
		/********** ?�?�t?�?�F?�?�b?�?�`?�?�f?�?�[?�?�^ **********/
		.inst		 (insn),				// ?�?�t?�?�F?�?�b?�?�`?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�
		/********** ?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�?�?�?�?�M?�?�?�?� **********/
		.stall		 (stall),				// ?�?�X?�?�g?�?�[?�?�?�?�
		.flush		 (flush),				// ?�?�t?�?�?�?�?�?�b?�?�V?�?�?�?�
		.new_pc		 (new_pc),				// ?�?�V?�?�?�?�?�?�?�?�?�?�v?�?�?�?�?�?�O?�?�?�?�?�?�?�?�?�?�J?�?�E?�?�?�?�?�?�^
		.br_taken	 (br_taken),			// ?�?�?�?�?�?�?�?�?�?�?�撰?�?�?�?�?�?�
		.br_addr	 (br_addr),				// ?�?�?�?�?�?�?�?�?�?�?�?�?�?�A?�?�h?�?�?�?�?�?�X
		/********** IF/ID?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�?�?�?�?�W?�?�X?�?�^ **********/
		.if_pc		 (if_pc),				// ?�?�v?�?�?�?�?�?�O?�?�?�?�?�?�?�?�?�?�J?�?�E?�?�?�?�?�?�^
		.if_inst	 (if_insn),				// ?�?�?�?�?�?�?�?�
		.if_en		 (if_en)				// ?�?�p?�?�C?�?�v?�?�?�?�?�?�C?�?�?�?�?�?�f?�?�[?�?�^?�?�?�朽?�?�?�
	);

endmodule
