`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/03/19 16:10:43
// Design Name:
// Module Name: IF_sim
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`define WORD 32  // 1word
`define WORD_ADDR_W 30  // address width 1word

`define GPR_ADDR_MSB 5-1

`define WORD_MSB `WORD-1
`define WORD_ADDR_MSB `WORD_ADDR_W-1
`define RegAddrBus `GPR_ADDR_MSB:0


module MEM_sim();
	reg				   clk=0;			// ????N????????????b????N
	reg				   reset;		// ???????????????????????????Z????b????g
  reg				   stall;		   // ???�X???�g???�[???�???�
	reg				   flush;		   // ???�t???�???�???�b???�V???�???�
	wire				   busy;		   // ???�r???�W???�[???�M???�???�
	/********** ???�t???�H???�???�???�[???�f???�B???�???�???�O **********/
	wire [`WORD_MSB:0] fwd_data;	   // ???�t???�H???�???�???�[???�f???�B???�???�???�O???�f???�[???�^
	/********** SPM???�C???�???�???�^???�t???�F???�[???�X **********/
	reg [`WORD_MSB:0] spm_rd_data;	   // ???�ǂݏo???�???�???�f???�[???�^
	wire [`WORD_ADDR_MSB:0] spm_addr;	   // ???�A???�h???�???�???�X
	wire				   spm_as_;		   // ???�A???�h???�???�???�X???�X???�g???�???�???�[???�u
	wire				   spm_rw;		   // ???�ǂ݁^???�???�???�???�
	wire [`WORD_MSB:0] spm_wr_data;	   // ???�???�???�???�???�???�???�݃f???�[???�^
	/********** ???�o???�X???�C???�???�???�^???�t???�F???�[???�X **********/
	reg [`WORD_MSB:0] bus_rd_data;	   // ???�ǂݏo???�???�???�f???�[???�^
	reg				   bus_rdy_;	   // ???�???�???�f???�B
	reg				   bus_grnt_;	   // ???�o???�X???�O???�???�???�???�???�g
	wire				   bus_req_;	   // ???�o???�X???�???�???�N???�G???�X???�g
	wire [`WORD_ADDR_MSB:0] bus_addr;	   // ???�A???�h???�???�???�X
	wire				   bus_as_;		   // ???�A???�h???�???�???�X???�X???�g???�???�???�[???�u
	wire				   bus_rw;		   // ???�ǂ݁^???�???�???�???�
	wire [`WORD_MSB:0] bus_wr_data;	   // ???�???�???�???�???�???�???�݃f???�[???�^
	/********** EX/MEM???�p???�C???�v???�???�???�C???�???�???�???�???�W???�X???�^ **********/
	reg [`WORD_ADDR_MSB:0] ex_pc;		   // ???�v???�???�???�O???�???�???�???�???�J???�E???�???�???�^
	reg				   ex_en;		   // ???�p???�C???�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
	reg				   ex_br_flag;	   // ???�???�???�???�???�t???�???�???�O
	reg [1:0]	   ex_mem_op;	   // ???�???�???�???�???�???�???�I???�y???�???�???�[???�V???�???�???�???�
	reg [`WORD_MSB:0] ex_mem_wr_data; // ???�???�???�???�???�???�???�???�???�???�???�???�???�݃f???�[???�^
	reg [1:0]   ex_ctrl_op;	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
	reg [4:0]  ex_dst_addr;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
	reg				   ex_gpr_we_;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
	reg [2:0]   ex_exp_code;	   // ???�???�???�O???�R???�[???�h
	reg [`WORD_MSB:0] ex_out;		   // ???�???�???�???�???�???�???�???�
	/********** MEM/WB???�p???�C???�v???�???�???�C???�???�???�???�???�W???�X???�^ **********/
	wire [`WORD_ADDR_MSB:0] mem_pc;		   // ???�v???�???�???�O???�???�???�???�???�J???�E???�???�???�^
	wire				   mem_en;		   // ???�p???�C???�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
	wire				   mem_br_flag;	   // ???�???�???�???�???�t???�???�???�O
	wire [1:0]   mem_ctrl_op;	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
	wire [4:0]  mem_dst_addr;   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
	wire				   mem_gpr_we_;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
	wire [2:0]   mem_exp_code;   // ???�???�???�O???�R???�[???�h
	wire [`WORD_MSB:0] mem_out;		   // ???�???�???�???�???�???�???�???�

    always begin
       clk=~clk; #(5);
    end
    stage_MEM stage_MEM (
    	/********** ???�N???�???�???�b???�N & ???�???�???�Z???�b???�g **********/
    	clk,			   // ???�N???�???�???�b???�N
    	reset,		   // ???�񓯊�???�???�???�Z???�b???�g
    	stall,		   // ???�X???�g???�[???�???�
    	flush,		   // ???�t???�???�???�b???�V???�???�
    	busy,		   // ???�r???�W???�[???�M???�???�
    	fwd_data,	   // ???�[???�f???�B???�???�???�O???�f???�[???�^
    	spm_rd_data,	   // ???�ǂݏo???�???�???�f???�[???�^
    	spm_addr,	   // ???�A???�h???�???�???�X
    	spm_as_,		   // ???�A???�h???�???�???�X???�X???�g???�???�???�[???�u
    	spm_rw,		   // ???�ǂ݁^???�???�???�???�
    	spm_wr_data,	   // ???�???�???�???�???�???�???�݃f???�[???�^
    	bus_rd_data,	   // ???�ǂݏo???�???�???�f???�[???�^
    	bus_rdy_,	   // ???�???�???�f???�B
    	bus_grnt_,	   // ???�o???�X???�O???�???�???�???�???�g
    	bus_req_,	   // ???�o???�X???�???�???�N???�G???�X???�g
    	bus_as_,		   // ???�A???�h???�???�???�X???�X???�g???�???�???�[???�u
    	bus_rw,		   // ???�ǂ݁^???�???�???�???�
    	bus_wr_data,	   // ???�???�???�???�???�???�???�݃f???�[???�^
    	ex_pc,		   // ???�???�???�???�???�J???�E???�???�???�^
    	ex_en,		   // �???�???�C???�???�???�f???�[???�^???�̗L???�???�
    	ex_br_flag,	   // ???�???�???�???�???�t???�???�???�O
    	ex_mem_op,	   // ?�???�???�I???�y???�???�???�[???�V???�???�???�???�
    	ex_mem_wr_data, // ?�???�???�???�???�???�???�???�???�݃f???�[???�^
    	ex_ctrl_op,	   // �X???�^???�I???�y???�???�???�[???�V???�???�???�???�
    	ex_dst_addr,	   // W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
    	ex_gpr_we_,	   // W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
    	ex_exp_code,	   // ???�???�???�O???�R???�[???�h
    	ex_out,		   // ???�???�???�???�???�???�???�???�
    	nem_pc,		   // ???�???�???�???�???�J???�E???�???�???�^
    	mem_en,		   // �???�???�C???�???�???�f???�[???�^???�̗L???�???�
    	mem_br_flag,	   // ???�???�???�???�???�t???�???�???�O
    	mem_ctrl_op,	   // �X???�^???�I???�y???�???�???�[???�V???�???�???�???�
    	mem_dst_addr,   // W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
    	mem_gpr_we_,	   // W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
    	mem_exp_code,   // ???�???�???�O???�R???�[???�h
    	mem_out		   // ???�???�???�???�???�???�???�???�
    );
  initial begin
    reset = 1;
		#(2)
    reset <= 0;
		repeat(2) @(posedge clk);
    reset <= 1;
		stall=0;
		flush=0;

    repeat(200) @(posedge clk);

    $stop;
  end

endmodule
