`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/03/19 16:10:43
// Design Name:
// Module Name: IF_sim
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`define WORD 32  // 1word
`define WORD_ADDR_W 30  // address width 1word

`define GPR_ADDR_MSB 5-1

`define WORD_MSB `WORD-1
`define WORD_ADDR_MSB `WORD_ADDR_W-1
`define RegAddrBus `GPR_ADDR_MSB:0


module EX_sim();
	reg				   clk=0;			// ????N????????????b????N
	reg				   reset;		// ???????????????????????????Z????b????g

  reg 				   stall;		   // ???�X???�g???�[???�???�
  reg 				   flush;		   // ???�t???�???�???�b???�V???�???�
  reg 				   int_detect;	   // ???�???�???�荞�݌�???�o
  reg  [`WORD_MSB:0] fwd_data;
  reg  [`WORD_ADDR_MSB:0] id_pc;		   // ???�v???�???�???�O???�???�???�???�???�J???�E???�???�???�^
  reg 				   id_en;		   // ???�p???�C???�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
  reg 				   id_br_flag;	   // ???�???�???�???�???�t???�???�???�O
  reg [3:0] id_alu_op;
  reg [`WORD_MSB:0] id_alu_in_0;
  reg [`WORD_MSB:0] id_alu_in_1;
  reg  [1:0]	   id_mem_op;	   // ???�???�???�???�???�???�???�I???�y???�???�???�[???�V???�???�???�???�
  reg  [`WORD_MSB:0] id_mem_wr_data; // ???�???�???�???�???�???�???�???�???�???�???�???�???�݃f???�[???�^
  reg  [1:0]   id_ctrl_op;	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
  reg  [`RegAddrBus]  id_dst_addr;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
  reg 				   id_gpr_we_;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
  reg  [2:0]   id_exp_code;	   // ???�???�???�O???�R???�[???�h
  /********** EX/MEM???�p???�C???�v???�???�???�C???�???�???�???�???�W???�X???�^ **********/
  wire [`WORD_ADDR_MSB:0] ex_pc;		   // ???�v???�???�???�O???�???�???�???�???�J???�E???�???�???�^
  wire				   ex_en;		   // ???�p???�C???�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
  wire				   ex_br_flag;	   // ???�???�???�???�???�t???�???�???�O
  wire [1:0]	   ex_mem_op;	   // ???�???�???�???�???�???�???�I???�y???�???�???�[???�V???�???�???�???�
  wire [`WORD_MSB:0] ex_mem_wr_data; // ???�???�???�???�???�???�???�???�???�???�???�???�???�݃f???�[???�^
  wire [1:0]   ex_ctrl_op;	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
  wire [`RegAddrBus]  ex_dst_addr;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�݃A???�h???�???�???�X
  wire				   ex_gpr_we_;	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
  wire [2:0]   ex_exp_code;	   // ???�???�???�O???�R???�[???�h
  wire [`WORD_MSB:0] ex_out;		   // ???�???�???�???�???�???�???�???�

  /********** ALU???�̏o???�???� **********/
  wire [`WORD_MSB:0]		   alu_out;		   // ???�???�???�Z???�???�???�???�
  wire					   alu_of;		   // ???�I???�[???�o???�t???�???�???�[

  /********** ???�???�???�Z???�???�???�ʂ̃t???�H???�???�???�[???�f???�B???�???�???�O **********/



  stage_EX ex(

	   clk,			   // ???�N???�???�???�b???�N
	   reset,		   // ???�񓯊�???�???�???�Z???�b???�g
	   stall,		   // ???�X???�g???�[???�???�
	   flush,		   // ???�t???�???�???�b???�V???�???�
	   int_detect,	   // ???�???�???�荞�݌�???�o
     fwd_data,
     id_pc,		   // ?�???�O???�???�???�???�???�J???�E???�???�???�^
	   id_en,		   // ??�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
	   id_br_flag,	   // ???�???�???�???�???�t???�???�???�O
     id_alu_op,
     id_alu_in_0,
     id_alu_in_1,
     id_mem_op,	   // �???�???�???�???�I???�y???�???�???�[???�V???�???�???�???�
     id_mem_wr_data, // �???�???�???�???�???�???�???�???�???�???�݃f???�[???�^
	id_ctrl_op,	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
	id_dst_addr,	   //    
	id_gpr_we_,	   // ???�ėp???�???�???�W???�X???�^???�???�???�???�???�???�???�ݗL???�???�
  	id_exp_code,	   // ???�???�???�O???�R???�[???�h
  	ex_pc,		   // ???�v???�???�???�O???�???�???�???�???�J???�E???�???�???�^
  	ex_en,		   // ???�p???�C???�v???�???�???�C???�???�???�f???�[???�^???�̗L???�???�
  	ex_br_flag,	   // ???�???�???�???�???�t???�???�???�O
  	ex_mem_op,	   // ???�???�???�???�???�???�???�I???�y???�???�???�[???�V???�???�???�???�
  	ex_mem_wr_data, // ???�???�???�???�???�???�???�???�???�???�???�???�???�݃f???�[???�^
  	ex_ctrl_op,	   // ???�???�???�䃌�W???�X???�^???�I???�y???�???�???�[???�V???�???�???�???�
  	ex_dst_addr,	   //
  	ex_gpr_we_,	   // ???�ėp???�???�???�W???�X???�???�
  	ex_exp_code,	   // ???�???�???�O???�R???�[???�h
  	ex_out		   // ???�???�???�???�???�???�???�???�
  );

    always begin
       clk=~clk; #(5);
    end


  initial begin
    reset = 1;
		#(2)
    reset <= 0;
		repeat(2) @(posedge clk);
    reset <= 1;
	 id_alu_in_0=10;
	 id_alu_in_1=20;
		stall=0;
		flush=0;
     repeat(200) @(posedge clk);
		stall=0;
		flush=1;
    repeat(200) @(posedge clk);
		stall=1;
		flush=0;
    repeat(200) @(posedge clk);
		stall=1;
		flush=1;
		repeat(200) @(posedge clk);
		stall=0;
		flush=0;
		repeat(200) @(posedge clk);

    repeat(200) @(posedge clk);

    $finish;
  end

endmodule
