`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/02/28 17:44:20
// Design Name: 
// Module Name: bus_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bus_sim(
    input clk,
    input rst,
    input mreq,
    input mgrnt,
    input mas,
    input mrw
    );
endmodule
