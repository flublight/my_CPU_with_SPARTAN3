`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/03/19 16:10:43
// Design Name:
// Module Name: IF_sim
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`define WORD 32  // 1word
`define WORD_ADDR_W 30  // address width 1word

`define GPR_ADDR_MSB 5-1

`define WORD_MSB `WORD-1
`define WORD_ADDR_MSB `WORD_ADDR_W-1
`define RegAddrBus `GPR_ADDR_MSB:0


module ID_sim();
	reg				   clk=0;			// ????N????????????b????N
	reg				   reset;		// ???????????????????????????Z????b????g

   reg [`WORD_MSB:0]	 gpr_rd_data_0;	 // ???o???f?[?^ 0
	reg [`WORD_MSB:0]	 gpr_rd_data_1;	 // ???o???f?[?^ 1
	wire [`GPR_ADDR_MSB:0]	 gpr_rd_addr_0;	 // ???o???A?h???X 0
	wire [`GPR_ADDR_MSB:0]	 gpr_rd_addr_1;	 // ???o???A?h???X 1
	/********** ?t?H???[?f?B???O **********/
	// EX?X?e?[?W??????t?H???[?f?B???O
	reg 					 ex_en;			// ?p?C?v???C???f?[?^??L??
	reg [`WORD_MSB:0]	 ex_fwd_data;	 // ?t?H???[?f?B???O?f?[?^
	reg [`GPR_ADDR_MSB:0]	 ex_dst_addr;	 // ????????A?h???X
	reg 					 ex_gpr_we_;	 // ????????L??
	// MEM?X?e?[?W??????t?H???[?f?B???O
	reg [`WORD_MSB:0]	 mem_fwd_data;	 // ?t?H???[?f?B???O?f?[?^
	/********** ?????W?X?^?C???^?t?F?[?X **********/
	reg exe_mode;		 // ???s???[?h
	reg [`WORD_MSB:0]	 creg_rd_data;	 // ???o???f?[?^
	wire [`GPR_ADDR_MSB:0]	 creg_rd_addr;	 // ???o???A?h???X
	/********** ?p?C?v???C???????M?? **********/
	reg 					 stall;			 // ?X?g?[??
	reg 					 flush;			 // ?t???b?V??
	wire [`WORD_ADDR_MSB:0]	 br_addr;		 // ?????A?h???X
	wire					 br_taken;		 // ?????????
	wire					 ld_hazard;		 // ???[?h?n?U?[?h
	/********** IF/ID?p?C?v???C?????W?X?^ **********/
	reg [`WORD_ADDR_MSB:0]	 if_pc;			 // ?v???O?????J?E???^
	reg [`WORD_MSB:0]	 if_insn;		 // ????
	reg 					 if_en;			 // ?p?C?v???C???f?[?^??L??
	/********** ID/EX?p?C?v???C?????W?X?^ **********/
	wire [`WORD_ADDR_MSB:0]	 id_pc;			 // ?v???O?????J?E???^
	wire					 id_en;			 // ?p?C?v???C???f?[?^??L??
	wire [3:0]		 id_alu_op;		 // ALU?I?y???[?V????
	wire [`WORD_MSB:0]	 id_alu_in_0;	 // ALU???? 0
	wire [`WORD_MSB:0]	 id_alu_in_1;	 // ALU???? 1
	wire					 id_br_flag;	 // ?????t???O
	wire [1:0]		 id_mem_op;		 // ???????I?y???[?V????
	wire [`WORD_MSB:0]	 id_mem_wr_data; // ??????????????f?[?^
	wire [1:0]	 id_ctrl_op;	 // ?????I?y???[?V????
	wire [`GPR_ADDR_MSB:0]	 id_dst_addr;	 // GPR????????A?h???X
	wire					 id_gpr_we_;	 // GPR????????L??
	wire [2:0]	 id_exp_code;	 // ???O?R?[?h


	/********** ?f?R?[?h?M?? **********/
	wire  [3:0]			 alu_op;		 // ALU?I?y???[?V????
	wire  [`WORD_MSB:0]		 alu_in_0;		 // ALU???? 0
	wire  [`WORD_MSB:0]		 alu_in_1;		 // ALU???? 1
	wire						 br_flag;		 // ?????t???O
	wire  [1:0]			 mem_op;		 // ???????I?y???[?V????
	wire  [`WORD_MSB:0]		 mem_wr_data;	 // ??????????????f?[?^
	wire  [1:0]			 ctrl_op;		 // ?????I?y???[?V????
	wire  [`GPR_ADDR_MSB:0]			 dst_addr;		 // GPR????????A?h???X
	wire						 gpr_we_;		 // GPR????????L??
	wire  [2:0]			 exp_code;		 // ???O?R?[?h

	stage_ID stage_ID(
 	 clk,			 // ?N???b?N
 	 reset,			 // ??????Z?b?g
 	 gpr_rd_data_0,	 // ???o???f?[?^ 0
 	 gpr_rd_data_1,	 // ???o???f?[?^ 1
 	 gpr_rd_addr_0,	 // ???o???A?h???X 0
 	 gpr_rd_addr_1,	 // ???o???A?h???X 1
 	 ex_en,			// ?p?C?v???C???f?[?^??L??
 	 ex_fwd_data,	 // ?t?H???[?f?B???O?f?[?^
 	 ex_dst_addr,	 // ????????A?h???X
 	 ex_gpr_we_,	 // ????????L??
 	 mem_fwd_data,	 // ?t?H???[?f?B???O?f?[?^
 	 exe_mode,		 // ???s???[?h
 	 creg_rd_data,	 // ???o???f?[?^
 	 creg_rd_addr,	 // ???o???A?h???X
	 stall,			 // ?X?g?[??
 	 flush,			 // ?t???b?V??
 	 br_addr,		 // ?????A?h???X
 	 br_taken,		 // ?????????
 	ld_hazard,		 // ???[?h?n?U?[?h
	 if_pc,			 // ?v???O?????J?E???^
 	 if_insn,		 // ????
 	 if_en,			 // ?p?C?v???C???f?[?^??L??
 	 id_pc,			 // ?v???O?????J?E???^
 	 id_en,			 // ?p?C?v???C???f?[?^??L??
 	 id_alu_op,		 // ALU?I?y???[?V????
 	 id_alu_in_0,	 // ALU???? 0
 	 id_alu_in_1,	 // ALU???? 1
 	 id_br_flag,	 // ?????t???O
 	 id_mem_op,		 // ???????I?y???[?V????
 	 id_mem_wr_data, // ??????????????f?[?^
 	 id_ctrl_op,	 // ?????I?y???[?V????
 	 id_dst_addr,	 // GPR????????A?h???X
 	 id_gpr_we_,	 // GPR????????L??
 	 id_exp_code	 // ???O?R?[?h
 );

    always begin
       clk=~clk; #(5);
    end


  initial begin
    reset = 1;
		#(2)
    reset <= 0;
		repeat(2) @(posedge clk);
    reset <= 1;
		stall=0;
  	flush=0;
    ex_en=1;
    ex_dst_addr=11;
    if_en=0;
    if_insn=3;
    if_pc=1000;
    repeat(200) @(posedge clk);
		stall=0;
		flush=1;
    repeat(200) @(posedge clk);
		stall=1;
		flush=0;
    repeat(200) @(posedge clk);
		stall=1;
		flush=1;
		repeat(200) @(posedge clk);
		stall=0;
		flush=0;
		repeat(200) @(posedge clk);

    repeat(200) @(posedge clk);

    $finish;
  end

endmodule
